/*
 * ECE385-HelperTools/PNG-To-Txt
 * Author: Rishi Thakkar
 *
 */

module  Wall_sprite
(
		input [1:0] data_In,
		input [7:0] write_address, read_address,
		input we, Clk,

		output logic [1:0] data_Out
);

// mem has width of 3 bits and a total of 225 addresses
logic [1:0] mem [0:224];

initial
begin
	 $readmemh("sprite_bytes/Wall.txt", mem);
end


always_ff @ (posedge Clk) begin
	if (we)
		mem[write_address] <= data_In;
	data_Out<= mem[read_address];
end

endmodule
