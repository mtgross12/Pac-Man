module Pac_valid_move(input next_x, next_y, sprite_num,
						output valid);
						
						